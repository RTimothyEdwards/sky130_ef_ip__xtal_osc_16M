magic
tech sky130A
magscale 1 2
timestamp 1699547177
<< dnwell >>
rect 116 112 9354 5580
<< nwell >>
rect 0 5374 9470 5696
rect 0 318 322 5374
rect 9148 318 9470 5374
rect 0 0 9470 318
<< psubdiff >>
rect 9978 5586 10902 5591
rect 9978 5548 10048 5586
rect 10835 5548 10902 5586
rect 9978 5541 10902 5548
rect 9978 5496 10028 5541
rect 9978 197 9987 5496
rect 10021 197 10028 5496
rect 9978 134 10028 197
rect 10852 5496 10902 5541
rect 10852 197 10861 5496
rect 10895 197 10902 5496
rect 10852 134 10902 197
rect 9978 128 10902 134
rect 9978 90 10055 128
rect 10842 90 10902 128
rect 9978 84 10902 90
<< mvnsubdiff >>
rect 73 5603 9397 5623
rect 73 5569 153 5603
rect 9317 5569 9397 5603
rect 73 5549 9397 5569
rect 73 5543 147 5549
rect 73 149 93 5543
rect 127 149 147 5543
rect 73 143 147 149
rect 9323 5543 9397 5549
rect 9323 149 9343 5543
rect 9377 149 9397 5543
rect 9323 143 9397 149
rect 73 123 9397 143
rect 73 89 153 123
rect 9317 89 9397 123
rect 73 69 9397 89
<< psubdiffcont >>
rect 10048 5548 10835 5586
rect 9987 197 10021 5496
rect 10861 197 10895 5496
rect 10055 90 10842 128
<< mvnsubdiffcont >>
rect 153 5569 9317 5603
rect 93 149 127 5543
rect 9343 149 9377 5543
rect 153 89 9317 123
<< locali >>
rect 93 5569 153 5603
rect 9317 5580 9575 5603
rect 9317 5569 9400 5580
rect 93 5554 233 5569
rect 93 5543 125 5554
rect 208 4045 233 5554
rect 9343 5543 9400 5569
rect 370 5422 7590 5440
rect 370 5366 410 5422
rect 2238 5416 7590 5422
rect 2238 5366 2574 5416
rect 7499 5366 7590 5416
rect 370 5302 7590 5366
rect 370 5295 4640 5302
rect 370 5292 2273 5295
rect 127 3301 233 4045
rect 203 2571 233 3301
rect 2184 2672 2273 5292
rect 2136 2668 2273 2672
rect 127 1577 233 2571
rect 372 2566 2273 2668
rect 2477 5292 4640 5295
rect 5085 5292 7590 5302
rect 2477 2672 2568 5292
rect 6839 4257 6978 5292
rect 6839 2680 6874 4257
rect 6941 2680 6978 4257
rect 2477 2668 2597 2672
rect 6839 2668 6978 2680
rect 7064 4684 7203 5292
rect 7064 2687 7097 4684
rect 7164 2687 7203 4684
rect 7064 2668 7203 2687
rect 2477 2664 4640 2668
rect 5085 2664 7207 2668
rect 2477 2566 7207 2664
rect 372 2526 7207 2566
rect 372 2457 1089 2526
rect 93 127 121 149
rect 202 127 233 1577
rect 839 2388 1089 2457
rect 839 422 913 2388
rect 1023 2269 1089 2388
rect 1549 2449 6404 2454
rect 1549 2444 4017 2449
rect 1549 2314 2834 2444
rect 3474 2319 4017 2444
rect 4657 2447 6404 2449
rect 4657 2319 5164 2447
rect 3474 2314 5164 2319
rect 1549 2311 5164 2314
rect 5563 2311 6404 2447
rect 1549 2300 6404 2311
rect 6498 2439 7207 2526
rect 1023 2156 1439 2269
rect 1023 1907 1089 2156
rect 1354 1907 1439 2156
rect 1023 1531 1439 1907
rect 1549 1850 1670 2300
rect 1549 1848 1958 1850
rect 1549 1700 1640 1848
rect 1780 1700 1958 1848
rect 2400 1848 6410 1850
rect 2400 1700 2704 1848
rect 1549 1699 2704 1700
rect 3618 1846 6410 1848
rect 3618 1699 3884 1846
rect 4239 1699 4505 1846
rect 4860 1699 6410 1846
rect 1549 1696 6410 1699
rect 1023 1530 1358 1531
rect 1023 422 1089 1530
rect 839 386 1089 422
rect 840 380 1089 386
rect 2085 1464 5946 1624
rect 2085 1034 2183 1464
rect 2085 1019 5948 1034
rect 2085 1018 5006 1019
rect 2085 880 2161 1018
rect 2308 880 2739 1018
rect 2886 1016 4375 1018
rect 2886 880 3300 1016
rect 2085 878 3300 880
rect 3447 880 4375 1016
rect 4522 881 5006 1018
rect 5829 881 5948 1019
rect 4522 880 5948 881
rect 3447 878 5948 880
rect 2085 874 5948 878
rect 2085 436 2183 874
rect 2085 417 5940 436
rect 2085 296 2162 417
rect 5912 296 5940 417
rect 2085 276 5940 296
rect 6498 413 6598 2439
rect 7050 2420 7207 2439
rect 7036 2335 7209 2420
rect 7036 1919 7041 2335
rect 7143 2263 7209 2335
rect 7485 2263 7586 5292
rect 7143 2117 7586 2263
rect 7143 1919 7209 2117
rect 7036 1261 7209 1919
rect 7035 1248 7308 1261
rect 7035 875 7045 1248
rect 7296 875 7308 1248
rect 7035 863 7308 875
rect 7036 566 7209 863
rect 7036 553 7515 566
rect 7036 413 7049 553
rect 6498 252 7049 413
rect 7036 218 7049 252
rect 7503 218 7515 553
rect 7036 204 7515 218
rect 93 123 233 127
rect 9377 149 9400 5543
rect 9343 123 9400 149
rect 93 89 153 123
rect 9317 117 9400 123
rect 9564 117 9575 5580
rect 9317 89 9575 117
rect 9801 5586 10902 5591
rect 9801 5572 10048 5586
rect 9801 125 9830 5572
rect 9962 5548 10048 5572
rect 10835 5548 10902 5586
rect 9962 5496 10902 5548
rect 9962 197 9987 5496
rect 10021 5477 10861 5496
rect 10021 5299 10120 5477
rect 10787 5299 10861 5477
rect 10021 4637 10861 5299
rect 10021 4171 10293 4637
rect 10021 2476 10028 4171
rect 10195 3310 10790 3326
rect 10195 3248 10498 3310
rect 10656 3248 10790 3310
rect 10195 3225 10790 3248
rect 10195 2907 10330 3225
rect 10852 2786 10861 4637
rect 10556 2764 10861 2786
rect 10021 2468 10207 2476
rect 10561 2468 10861 2764
rect 10021 2452 10861 2468
rect 10021 2403 10055 2452
rect 10413 2403 10861 2452
rect 10021 2362 10861 2403
rect 10021 1522 10028 2362
rect 10021 1030 10308 1522
rect 10852 1030 10861 2362
rect 10021 364 10861 1030
rect 10021 197 10111 364
rect 9962 186 10111 197
rect 10679 197 10861 364
rect 10895 197 10902 5496
rect 10679 186 10902 197
rect 9962 128 10902 186
rect 9962 125 10055 128
rect 9801 90 10055 125
rect 10842 90 10902 128
rect 9801 84 10902 90
<< viali >>
rect 125 5543 208 5554
rect 125 4045 127 5543
rect 127 4045 208 5543
rect 410 5366 2238 5422
rect 2574 5366 7499 5416
rect 121 2571 127 3301
rect 127 2571 203 3301
rect 2273 2566 2477 5295
rect 6874 2680 6941 4257
rect 7097 2687 7164 4684
rect 121 149 127 1577
rect 127 149 202 1577
rect 121 127 202 149
rect 913 422 1023 2388
rect 2834 2314 3474 2444
rect 4017 2319 4657 2449
rect 5164 2311 5563 2447
rect 1640 1700 1780 1848
rect 1958 1700 2400 1850
rect 2704 1699 3618 1848
rect 3884 1699 4239 1846
rect 4505 1699 4860 1846
rect 2161 880 2308 1018
rect 2739 880 2886 1018
rect 3300 878 3447 1016
rect 4375 880 4522 1018
rect 5006 881 5829 1019
rect 2162 296 5912 417
rect 7041 1919 7143 2335
rect 7045 875 7296 1248
rect 7049 218 7503 553
rect 9400 117 9564 5580
rect 9830 125 9962 5572
rect 10120 5299 10787 5477
rect 10498 3248 10656 3310
rect 10055 2403 10413 2452
rect 10111 186 10679 364
<< metal1 >>
rect 119 5554 214 5566
rect 115 4045 125 5554
rect 208 4045 218 5554
rect 341 5422 9148 5439
rect 341 5366 410 5422
rect 2238 5416 9148 5422
rect 2238 5366 2574 5416
rect 7499 5366 9148 5416
rect 341 5295 9148 5366
rect 341 5294 2273 5295
rect 504 4768 740 5200
rect 836 4768 1072 5200
rect 1168 4768 1404 5200
rect 1500 4768 1736 5200
rect 1832 4768 2068 5200
rect 119 4033 214 4045
rect 0 3568 200 3656
rect 0 3533 314 3568
rect 0 3456 200 3533
rect 109 3301 220 3322
rect 109 2571 121 3301
rect 203 2571 220 3301
rect 109 2554 220 2571
rect 279 2507 314 3533
rect 378 3186 574 3200
rect 378 2785 392 3186
rect 555 2785 574 3186
rect 378 2768 574 2785
rect 670 2768 906 3200
rect 1002 2768 1238 3200
rect 1334 2768 1570 3200
rect 1666 2768 1902 3200
rect 2012 2824 2049 2842
rect 2012 2769 2060 2824
rect 636 2579 646 2644
rect 847 2579 857 2644
rect 261 2442 271 2507
rect 472 2442 482 2507
rect 676 2319 719 2579
rect 2012 2562 2049 2769
rect 1487 2525 2049 2562
rect 2234 2566 2273 5294
rect 2477 5294 9148 5295
rect 2477 2566 2523 5294
rect 2674 4767 2910 5199
rect 3006 4767 3242 5199
rect 3338 4767 3574 5199
rect 3670 4767 3906 5199
rect 4002 4767 4238 5199
rect 4334 4767 4570 5199
rect 4666 4767 4902 5199
rect 4998 4767 5234 5199
rect 5330 4767 5566 5199
rect 5662 4767 5898 5199
rect 5994 4767 6230 5199
rect 6326 4767 6562 5199
rect 6658 4833 6728 5199
rect 6968 5193 7377 5199
rect 6658 4789 6933 4833
rect 6658 4766 6728 4789
rect 6889 4544 6933 4789
rect 6968 4770 6992 5193
rect 7164 4770 7377 5193
rect 6968 4766 7377 4770
rect 7091 4695 7170 4696
rect 7082 4684 7178 4695
rect 6869 4338 6879 4544
rect 6937 4338 6947 4544
rect 6860 4257 6956 4272
rect 2674 3135 2722 3185
rect 2681 2767 2735 2843
rect 2840 2767 3076 3199
rect 3172 2767 3408 3199
rect 3504 2767 3740 3199
rect 3836 2767 4072 3199
rect 4168 2767 4404 3199
rect 4500 2767 4736 3199
rect 4832 2767 5068 3199
rect 5164 2767 5400 3199
rect 5496 2767 5732 3199
rect 5828 2767 6064 3199
rect 6160 2767 6396 3199
rect 6492 2767 6728 3199
rect 2234 2545 2523 2566
rect 1103 2444 1113 2509
rect 1314 2444 1324 2509
rect 898 2388 1033 2402
rect 0 1861 200 1918
rect 0 1800 414 1861
rect 0 1718 200 1800
rect 106 1577 218 1594
rect 106 127 121 1577
rect 202 127 218 1577
rect 353 933 414 1800
rect 353 872 728 933
rect 898 422 913 2388
rect 1023 422 1033 2388
rect 1197 1773 1244 2444
rect 1197 1726 1381 1773
rect 1334 1243 1381 1726
rect 1487 1273 1524 2525
rect 2687 2496 2725 2767
rect 6658 2766 6728 2767
rect 6860 2680 6874 4257
rect 6941 2680 6956 4257
rect 4723 2670 5169 2671
rect 2818 2668 3994 2669
rect 4723 2668 5571 2670
rect 2818 2661 5571 2668
rect 6860 2664 6956 2680
rect 7082 2687 7097 4684
rect 7164 2687 7178 4684
rect 9259 4642 9284 5609
rect 9595 4642 9617 5609
rect 7082 2667 7178 2687
rect 7580 3782 7702 3818
rect 2818 2654 4991 2661
rect 2818 2555 3985 2654
rect 2527 2431 2537 2496
rect 2738 2431 2748 2496
rect 2818 2444 3487 2555
rect 2818 2314 2834 2444
rect 3474 2314 3487 2444
rect 3534 2443 3544 2508
rect 3745 2443 3755 2508
rect 2818 2313 3487 2314
rect 2822 2308 3486 2313
rect 1703 1860 1784 2117
rect 1634 1848 1786 1860
rect 1630 1700 1640 1848
rect 1780 1700 1790 1848
rect 1634 1688 1786 1700
rect 1847 1391 1883 2202
rect 1944 2168 3145 2206
rect 1944 2028 1982 2168
rect 2321 1856 2402 2117
rect 2466 1961 2498 2168
rect 1946 1850 2412 1856
rect 1946 1700 1958 1850
rect 2400 1700 2412 1850
rect 1946 1694 2412 1700
rect 2572 1531 2618 2168
rect 2937 1854 3018 2115
rect 3077 1960 3109 2168
rect 3181 2055 3635 2091
rect 2692 1848 3630 1854
rect 2692 1699 2704 1848
rect 3618 1699 3630 1848
rect 2692 1693 3630 1699
rect 2572 1485 3066 1531
rect 3703 1507 3738 2443
rect 3964 2401 3985 2555
rect 4769 2409 4991 2654
rect 5551 2453 5571 2661
rect 5784 2552 5794 2617
rect 5995 2552 6005 2617
rect 6055 2563 7329 2597
rect 5551 2447 5575 2453
rect 4769 2401 5164 2409
rect 3964 2319 4017 2401
rect 4657 2366 5164 2401
rect 4657 2319 4790 2366
rect 3964 2313 4790 2319
rect 3964 2119 4240 2313
rect 3797 1569 3839 2117
rect 3964 1852 4241 2119
rect 3872 1846 4251 1852
rect 3872 1699 3884 1846
rect 4239 1699 4251 1846
rect 3872 1693 4251 1699
rect 4316 1569 4353 2192
rect 4526 2121 4790 2313
rect 4875 2249 4885 2314
rect 5086 2249 5096 2314
rect 5144 2311 5164 2366
rect 5563 2311 5575 2447
rect 5705 2433 5715 2462
rect 5144 2305 5575 2311
rect 5654 2397 5715 2433
rect 5916 2397 5926 2462
rect 5144 2304 5571 2305
rect 4409 1663 4446 2117
rect 4526 1852 4866 2121
rect 4493 1846 4872 1852
rect 4493 1699 4505 1846
rect 4860 1699 4872 1846
rect 4493 1693 4872 1699
rect 4409 1658 4727 1663
rect 4935 1658 4971 2187
rect 5035 1784 5075 2249
rect 5253 2028 5263 2121
rect 5505 2028 5515 2121
rect 5035 1744 5285 1784
rect 4409 1626 5176 1658
rect 4690 1622 5176 1626
rect 3797 1532 4624 1569
rect 3530 1486 3540 1507
rect 1777 1326 1787 1391
rect 1988 1326 1998 1391
rect 2542 1368 2552 1385
rect 2357 1332 2552 1368
rect 1487 1236 2307 1273
rect 2360 1150 2398 1332
rect 2542 1320 2552 1332
rect 2753 1368 2763 1385
rect 2753 1332 2950 1368
rect 2753 1320 2763 1332
rect 2149 1018 2320 1024
rect 2149 880 2161 1018
rect 2308 880 2320 1018
rect 2149 874 2320 880
rect 2236 608 2296 874
rect 2358 542 2394 742
rect 2464 542 2508 1300
rect 2808 1098 2852 1298
rect 2912 1144 2950 1332
rect 3020 1210 3066 1485
rect 3474 1442 3540 1486
rect 3741 1442 3751 1507
rect 3362 1100 3406 1294
rect 3474 1138 3509 1442
rect 3797 1288 3839 1532
rect 3571 1246 3840 1288
rect 3571 1205 3613 1246
rect 2808 1054 3068 1098
rect 3362 1056 3622 1100
rect 2727 1018 2898 1024
rect 2727 880 2739 1018
rect 2886 880 2898 1018
rect 2727 874 2898 880
rect 2784 610 2844 874
rect 2918 542 2954 748
rect 3024 608 3068 1054
rect 3288 1016 3459 1022
rect 3288 878 3300 1016
rect 3447 878 3459 1016
rect 3288 872 3459 878
rect 3348 608 3408 872
rect 3474 546 3510 754
rect 3578 606 3622 1056
rect 4447 1024 4524 1294
rect 4587 1166 4624 1532
rect 4690 1205 4727 1622
rect 4806 1437 4816 1502
rect 5017 1437 5027 1502
rect 4363 1018 4534 1024
rect 4363 880 4375 1018
rect 4522 880 4534 1018
rect 4582 970 4625 1166
rect 4582 927 4734 970
rect 4363 874 4534 880
rect 4447 870 4524 874
rect 4032 784 4066 786
rect 4220 784 4230 797
rect 4024 746 4230 784
rect 3753 629 3975 669
rect 3753 542 3793 629
rect 4032 547 4066 746
rect 4220 732 4230 746
rect 4431 784 4441 797
rect 4431 746 4648 784
rect 4431 732 4441 746
rect 2336 502 3793 542
rect 4133 435 4205 698
rect 4440 435 4523 690
rect 4585 544 4619 746
rect 4691 603 4734 927
rect 4875 668 4915 1437
rect 5006 1025 5083 1298
rect 5140 1163 5176 1622
rect 5245 1207 5285 1744
rect 5545 1655 5577 2182
rect 5654 1749 5690 2397
rect 5954 2059 5986 2552
rect 5904 2027 5986 2059
rect 6055 2029 6089 2563
rect 6156 2457 7254 2493
rect 5654 1713 5835 1749
rect 5545 1623 5730 1655
rect 5698 1376 5730 1623
rect 5400 1340 5731 1376
rect 5400 1163 5436 1340
rect 5140 1127 5436 1163
rect 5550 1025 5627 1299
rect 5698 1142 5730 1340
rect 5799 1204 5835 1713
rect 4994 1019 5841 1025
rect 4994 881 5006 1019
rect 5829 881 5841 1019
rect 4994 875 5841 881
rect 5006 874 5083 875
rect 5122 794 5764 798
rect 5904 794 5936 2027
rect 6156 1976 6192 2457
rect 7035 2342 7149 2347
rect 6869 2335 7150 2342
rect 6277 2104 6719 2117
rect 6256 2052 6726 2104
rect 6277 2049 6719 2052
rect 6011 1880 6051 1889
rect 6004 1815 6014 1880
rect 6215 1815 6225 1880
rect 5122 762 5936 794
rect 5122 754 5764 762
rect 4875 628 5091 668
rect 5136 533 5174 752
rect 5247 503 5330 691
rect 5552 503 5635 689
rect 5697 542 5735 754
rect 6011 671 6051 1815
rect 6277 1728 6345 2049
rect 6869 1919 7041 2335
rect 7143 1919 7150 2335
rect 7218 2302 7254 2457
rect 7580 2302 7616 3782
rect 7644 3563 7654 3628
rect 7855 3563 7865 3628
rect 9259 3077 9400 4642
rect 9137 2400 9400 3077
rect 7218 2266 7616 2302
rect 7646 2068 7656 2133
rect 7857 2068 7867 2133
rect 6869 1909 7150 1919
rect 7035 1907 7149 1909
rect 7646 1841 7656 1906
rect 7857 1841 7867 1906
rect 5784 631 6051 671
rect 6094 1660 6345 1728
rect 5247 502 5635 503
rect 6094 502 6162 1660
rect 7035 1248 7308 1261
rect 6703 509 6939 941
rect 7035 875 7045 1248
rect 7296 875 7308 1248
rect 7035 863 7308 875
rect 7036 554 9224 566
rect 7036 553 7897 554
rect 5247 464 6162 502
rect 5247 435 5330 436
rect 5552 435 5635 436
rect 898 408 1033 422
rect 2138 417 5941 435
rect 2138 296 2162 417
rect 5912 296 5941 417
rect 2138 276 5941 296
rect 7036 218 7049 553
rect 7503 218 7897 553
rect 7036 216 7897 218
rect 9111 216 9224 554
rect 7036 204 9224 216
rect 106 109 218 127
rect 9259 117 9400 2400
rect 9564 117 9617 4642
rect 9259 84 9617 117
rect 9780 5572 10902 5596
rect 9780 125 9830 5572
rect 9962 5477 10902 5572
rect 9962 5299 10120 5477
rect 10787 5299 10902 5477
rect 9962 4636 10902 5299
rect 9962 2541 10085 4636
rect 10704 4014 10904 4214
rect 10252 3623 10904 3630
rect 10252 3439 10264 3623
rect 10723 3439 10904 3623
rect 10252 3430 10904 3439
rect 10479 3310 10682 3430
rect 10479 3248 10498 3310
rect 10656 3248 10682 3310
rect 10479 3134 10682 3248
rect 10386 2951 10425 3115
rect 10310 2912 10425 2951
rect 10310 2867 10349 2912
rect 10139 2802 10149 2867
rect 10350 2802 10360 2867
rect 10510 2853 10554 3055
rect 10443 2809 10554 2853
rect 10310 2599 10349 2802
rect 10443 2708 10487 2809
rect 10704 2708 10904 2728
rect 10443 2641 10904 2708
rect 10443 2640 10487 2641
rect 10381 2544 10497 2562
rect 10380 2541 10497 2544
rect 9962 2452 10499 2541
rect 10704 2528 10904 2641
rect 9962 2403 10055 2452
rect 10413 2403 10499 2452
rect 9962 2357 10499 2403
rect 9962 1056 10085 2357
rect 10255 2245 10737 2261
rect 10255 2078 10273 2245
rect 10721 2078 10737 2245
rect 10255 2063 10737 2078
rect 10704 1478 10904 1678
rect 9962 364 10904 1056
rect 9962 186 10111 364
rect 10679 186 10904 364
rect 9962 125 10904 186
rect 9780 92 10904 125
rect 9780 91 10085 92
<< via1 >>
rect 125 4045 208 5554
rect 392 2785 555 3186
rect 646 2579 847 2644
rect 271 2442 472 2507
rect 6992 4770 7164 5193
rect 6879 4338 6937 4544
rect 1113 2444 1314 2509
rect 913 422 1021 1635
rect 9284 5580 9595 5609
rect 9284 4642 9400 5580
rect 9400 4642 9564 5580
rect 9564 4642 9595 5580
rect 2537 2431 2738 2496
rect 3544 2443 3745 2508
rect 1640 1700 1780 1848
rect 1958 1700 2400 1850
rect 2704 1699 3618 1848
rect 3985 2449 4769 2654
rect 3985 2401 4017 2449
rect 4017 2401 4657 2449
rect 4657 2401 4769 2449
rect 4991 2447 5551 2661
rect 5794 2552 5995 2617
rect 4991 2409 5164 2447
rect 5164 2409 5551 2447
rect 3884 1699 4239 1846
rect 4885 2249 5086 2314
rect 5715 2397 5916 2462
rect 4505 1699 4860 1846
rect 5263 2028 5505 2121
rect 1787 1326 1988 1391
rect 2552 1320 2753 1385
rect 2161 880 2308 1018
rect 3540 1442 3741 1507
rect 2739 880 2886 1018
rect 3300 878 3447 1016
rect 4816 1437 5017 1502
rect 4375 880 4522 1018
rect 4230 732 4431 797
rect 5006 881 5829 1019
rect 6014 1815 6215 1880
rect 7654 3563 7855 3628
rect 7656 2068 7857 2133
rect 7656 1841 7857 1906
rect 7045 875 7296 1248
rect 2162 296 5912 417
rect 7049 218 7503 553
rect 7897 216 9111 554
rect 10264 3439 10723 3623
rect 10149 2802 10350 2867
rect 10273 2078 10721 2245
<< metal2 >>
rect 7469 5655 9615 5657
rect 0 5609 9615 5655
rect 0 5554 9284 5609
rect 0 4045 125 5554
rect 208 5193 9284 5554
rect 208 4770 6992 5193
rect 7164 4770 9284 5193
rect 208 4642 9284 4770
rect 9595 4642 9615 5609
rect 208 4617 9615 4642
rect 208 4045 6681 4617
rect 6879 4544 6937 4554
rect 6879 4328 6937 4338
rect 0 4027 6681 4045
rect 342 3186 596 4027
rect 342 2785 392 3186
rect 555 2785 596 3186
rect 342 2734 596 2785
rect 3966 3653 4796 4027
rect 4960 3653 5573 4027
rect 3966 2654 4794 3653
rect 646 2644 847 2654
rect 847 2591 3856 2631
rect 646 2569 847 2579
rect 271 2507 472 2517
rect 1113 2509 1314 2519
rect 472 2457 1113 2492
rect 271 2432 472 2442
rect 3544 2508 3745 2518
rect 2537 2496 2738 2506
rect 1314 2457 2537 2492
rect 1113 2434 1314 2444
rect 2738 2457 3544 2492
rect 3544 2433 3745 2443
rect 2537 2421 2738 2431
rect 3816 2301 3856 2591
rect 3966 2401 3985 2654
rect 4769 2401 4794 2654
rect 3966 2384 4794 2401
rect 4962 2661 5573 3653
rect 6886 2735 6926 4328
rect 7654 3628 7855 3638
rect 4962 2409 4991 2661
rect 5551 2409 5573 2661
rect 4962 2390 5573 2409
rect 5634 2695 6926 2735
rect 7394 3565 7654 3615
rect 4885 2314 5086 2324
rect 3816 2261 4885 2301
rect 5634 2301 5674 2695
rect 5794 2627 5839 2628
rect 5794 2624 5995 2627
rect 7394 2624 7444 3565
rect 10252 3623 10904 3630
rect 7855 3565 7918 3615
rect 7654 3553 7855 3563
rect 10252 3439 10264 3623
rect 10723 3439 10904 3623
rect 10252 3430 10904 3439
rect 10149 2867 10350 2877
rect 5794 2617 7444 2624
rect 5995 2574 7444 2617
rect 7497 2813 10149 2857
rect 5794 2542 5995 2552
rect 7497 2492 7541 2813
rect 10149 2792 10350 2802
rect 10428 2858 10904 3430
rect 5715 2462 5916 2472
rect 6212 2452 7541 2492
rect 5916 2448 7541 2452
rect 5916 2408 6256 2448
rect 5715 2387 5916 2397
rect 10428 2386 10736 2858
rect 5086 2261 6060 2301
rect 4885 2239 5086 2249
rect 5263 2121 5509 2131
rect 5505 2028 5509 2121
rect 1503 1850 4899 1972
rect 1503 1848 1958 1850
rect 1503 1700 1640 1848
rect 1780 1700 1958 1848
rect 2400 1848 4899 1850
rect 2400 1700 2704 1848
rect 1503 1699 2704 1700
rect 3618 1846 4899 1848
rect 3618 1699 3884 1846
rect 4239 1699 4505 1846
rect 4860 1699 4899 1846
rect 0 1635 1283 1650
rect 0 422 913 1635
rect 1021 1260 1283 1635
rect 1503 1601 4899 1699
rect 5263 1741 5509 2028
rect 6020 1890 6060 2261
rect 6330 2261 10736 2386
rect 6330 2245 10737 2261
rect 6330 2231 10273 2245
rect 6014 1880 6215 1890
rect 6014 1805 6215 1815
rect 6330 1741 6526 2231
rect 7656 2133 7857 2143
rect 5263 1578 6526 1741
rect 7235 2077 7656 2127
rect 3540 1507 3741 1517
rect 4816 1502 5017 1512
rect 3741 1451 4816 1486
rect 3540 1432 3741 1442
rect 4816 1427 5017 1437
rect 1787 1391 1988 1401
rect 2552 1385 2753 1395
rect 1988 1331 2552 1381
rect 1787 1316 1988 1326
rect 7235 1381 7285 2077
rect 7857 2077 7909 2127
rect 10255 2078 10273 2231
rect 10721 2078 10737 2245
rect 7656 2058 7857 2068
rect 10255 2063 10737 2078
rect 7656 1906 7857 1916
rect 2753 1331 7285 1381
rect 7359 1854 7656 1904
rect 2552 1310 2753 1320
rect 7035 1260 7308 1261
rect 1021 1248 7308 1260
rect 1021 1019 7045 1248
rect 1021 1018 5006 1019
rect 1021 880 2161 1018
rect 2308 880 2739 1018
rect 2886 1016 4375 1018
rect 2886 880 3300 1016
rect 1021 878 3300 880
rect 3447 880 4375 1016
rect 4522 881 5006 1018
rect 5829 881 7045 1019
rect 4522 880 7045 881
rect 3447 878 7045 880
rect 1021 875 7045 878
rect 7296 875 7308 1248
rect 1021 863 7308 875
rect 1021 862 7255 863
rect 1021 566 1654 862
rect 4230 797 4431 807
rect 7359 790 7409 1854
rect 7857 1854 7915 1904
rect 7656 1831 7857 1841
rect 4431 740 7409 790
rect 4230 722 4431 732
rect 1021 554 9222 566
rect 1021 553 7897 554
rect 1021 422 7049 553
rect 0 417 7049 422
rect 0 296 2162 417
rect 5912 296 7049 417
rect 0 218 7049 296
rect 7503 218 7897 553
rect 0 216 7897 218
rect 9111 216 9222 554
rect 0 25 9222 216
use sky130_fd_pr__diode_pd2nw_05v5_K4SERG  D1
timestamp 1698886478
transform 1 0 1357 0 1 1263
box -321 -321 321 321
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D2
timestamp 1698886478
transform 1 0 1219 0 1 2030
box -183 -183 183 183
use level_shifter  level_shifter_0
timestamp 1698887706
transform -1 0 10312 0 1 2782
box -422 -2464 2656 76
use level_shifter  level_shifter_1
timestamp 1698887706
transform -1 0 10312 0 -1 2910
box -422 -2464 2656 76
use sky130_fd_pr__pfet_01v8_LGS3BL  sky130_fd_pr__pfet_01v8_LGS3BL_0
timestamp 1698716925
transform 0 1 10542 -1 0 3083
box -211 -284 211 284
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM1
timestamp 1698886478
transform 1 0 3490 0 1 1250
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM2
timestamp 1698886478
transform 1 0 3714 0 1 2073
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM3
timestamp 1698886478
transform 1 0 4330 0 1 2073
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM4
timestamp 1698886478
transform 1 0 4602 0 1 1250
box -278 -300 278 300
use sky130_fd_pr__nfet_01v8_L9WNCD  XM5
timestamp 1699029959
transform 0 1 10399 -1 0 2609
box -211 -229 211 229
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM9
timestamp 1698886478
transform 1 0 4946 0 1 2073
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM10
timestamp 1698886478
transform 1 0 5158 0 1 1250
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM11
timestamp 1698886478
transform 1 0 5562 0 1 2073
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM12
timestamp 1698886478
transform 1 0 5714 0 1 1250
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM13
timestamp 1698886478
transform 1 0 4602 0 1 650
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM14
timestamp 1698886478
transform 1 0 6178 0 1 2073
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM21
timestamp 1698886478
transform 1 0 2378 0 1 650
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM22
timestamp 1698886478
transform 1 0 2482 0 1 2073
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM23
timestamp 1698886478
transform 1 0 2378 0 1 1250
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM24
timestamp 1698886478
transform 1 0 3098 0 1 2073
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM29
timestamp 1698886478
transform 1 0 3490 0 1 650
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM30
timestamp 1698886478
transform 1 0 2934 0 1 650
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM31
timestamp 1698886478
transform 1 0 5158 0 1 650
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM33
timestamp 1698886478
transform 1 0 4046 0 1 650
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM34
timestamp 1698886478
transform 1 0 1866 0 1 2073
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM36
timestamp 1698886478
transform 1 0 2934 0 1 1250
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM39
timestamp 1698886478
transform 1 0 5714 0 1 650
box -278 -300 278 300
use sky130_fd_pr__res_xhigh_po_0p35_CWLS5Y  XR1
timestamp 1698886478
transform 1 0 1286 0 1 3984
box -948 -1382 948 1382
use sky130_fd_pr__res_xhigh_po_0p35_7RFGLT  XR2
timestamp 1698886478
transform 1 0 696 0 1 1428
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_4FEQLC  XR3
timestamp 1698886478
transform 1 0 4701 0 1 3982
box -2193 -1382 2193 1382
use sky130_fd_pr__res_xhigh_po_0p35_ENTFM9  XR4
timestamp 1699029959
transform 1 0 6821 0 1 1425
box -284 -1082 284 1082
use sky130_fd_pr__res_xhigh_po_0p35_KNBXRF  XR5
timestamp 1698886478
transform 1 0 7341 0 1 3782
box -201 -1582 201 1582
<< labels >>
flabel metal2 0 25 202 1650 0 FreeSans 256 0 0 0 avss
port 3 nsew
flabel metal1 0 1718 200 1918 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 0 3456 200 3656 0 FreeSans 256 0 0 0 in
port 0 nsew
flabel metal2 0 4027 125 5655 0 FreeSans 256 0 0 0 avdd
port 2 nsew
flabel metal2 10726 2858 10904 3630 0 FreeSans 256 0 0 0 dvdd
port 4 nsew
flabel metal1 10708 92 10904 1056 0 FreeSans 256 0 0 0 dvss
port 5 nsew
flabel metal1 10704 1478 10904 1678 0 FreeSans 256 0 0 0 ena
port 6 nsew
flabel metal1 10704 4014 10904 4214 0 FreeSans 256 0 0 0 stdby
port 8 nsew
flabel metal1 10704 2528 10904 2728 0 FreeSans 256 0 0 0 dout
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 10904 5696
<< end >>
