magic
tech sky130A
magscale 1 2
timestamp 1698886478
<< pwell >>
rect -2193 -1382 2193 1382
<< psubdiff >>
rect -2157 1312 -2061 1346
rect 2061 1312 2157 1346
rect -2157 1250 -2123 1312
rect 2123 1250 2157 1312
rect -2157 -1312 -2123 -1250
rect 2123 -1312 2157 -1250
rect -2157 -1346 -2061 -1312
rect 2061 -1346 2157 -1312
<< psubdiffcont >>
rect -2061 1312 2061 1346
rect -2157 -1250 -2123 1250
rect 2123 -1250 2157 1250
rect -2061 -1346 2061 -1312
<< xpolycontact >>
rect -2027 784 -1957 1216
rect -2027 -1216 -1957 -784
rect -1861 784 -1791 1216
rect -1861 -1216 -1791 -784
rect -1695 784 -1625 1216
rect -1695 -1216 -1625 -784
rect -1529 784 -1459 1216
rect -1529 -1216 -1459 -784
rect -1363 784 -1293 1216
rect -1363 -1216 -1293 -784
rect -1197 784 -1127 1216
rect -1197 -1216 -1127 -784
rect -1031 784 -961 1216
rect -1031 -1216 -961 -784
rect -865 784 -795 1216
rect -865 -1216 -795 -784
rect -699 784 -629 1216
rect -699 -1216 -629 -784
rect -533 784 -463 1216
rect -533 -1216 -463 -784
rect -367 784 -297 1216
rect -367 -1216 -297 -784
rect -201 784 -131 1216
rect -201 -1216 -131 -784
rect -35 784 35 1216
rect -35 -1216 35 -784
rect 131 784 201 1216
rect 131 -1216 201 -784
rect 297 784 367 1216
rect 297 -1216 367 -784
rect 463 784 533 1216
rect 463 -1216 533 -784
rect 629 784 699 1216
rect 629 -1216 699 -784
rect 795 784 865 1216
rect 795 -1216 865 -784
rect 961 784 1031 1216
rect 961 -1216 1031 -784
rect 1127 784 1197 1216
rect 1127 -1216 1197 -784
rect 1293 784 1363 1216
rect 1293 -1216 1363 -784
rect 1459 784 1529 1216
rect 1459 -1216 1529 -784
rect 1625 784 1695 1216
rect 1625 -1216 1695 -784
rect 1791 784 1861 1216
rect 1791 -1216 1861 -784
rect 1957 784 2027 1216
rect 1957 -1216 2027 -784
<< xpolyres >>
rect -2027 -784 -1957 784
rect -1861 -784 -1791 784
rect -1695 -784 -1625 784
rect -1529 -784 -1459 784
rect -1363 -784 -1293 784
rect -1197 -784 -1127 784
rect -1031 -784 -961 784
rect -865 -784 -795 784
rect -699 -784 -629 784
rect -533 -784 -463 784
rect -367 -784 -297 784
rect -201 -784 -131 784
rect -35 -784 35 784
rect 131 -784 201 784
rect 297 -784 367 784
rect 463 -784 533 784
rect 629 -784 699 784
rect 795 -784 865 784
rect 961 -784 1031 784
rect 1127 -784 1197 784
rect 1293 -784 1363 784
rect 1459 -784 1529 784
rect 1625 -784 1695 784
rect 1791 -784 1861 784
rect 1957 -784 2027 784
<< locali >>
rect -2157 1312 -2061 1346
rect 2061 1312 2157 1346
rect -2157 1250 -2123 1312
rect 2123 1250 2157 1312
rect -2157 -1312 -2123 -1250
rect 2123 -1312 2157 -1250
rect -2157 -1346 -2061 -1312
rect 2061 -1346 2157 -1312
<< viali >>
rect -2011 801 -1973 1198
rect -1845 801 -1807 1198
rect -1679 801 -1641 1198
rect -1513 801 -1475 1198
rect -1347 801 -1309 1198
rect -1181 801 -1143 1198
rect -1015 801 -977 1198
rect -849 801 -811 1198
rect -683 801 -645 1198
rect -517 801 -479 1198
rect -351 801 -313 1198
rect -185 801 -147 1198
rect -19 801 19 1198
rect 147 801 185 1198
rect 313 801 351 1198
rect 479 801 517 1198
rect 645 801 683 1198
rect 811 801 849 1198
rect 977 801 1015 1198
rect 1143 801 1181 1198
rect 1309 801 1347 1198
rect 1475 801 1513 1198
rect 1641 801 1679 1198
rect 1807 801 1845 1198
rect 1973 801 2011 1198
rect -2011 -1198 -1973 -801
rect -1845 -1198 -1807 -801
rect -1679 -1198 -1641 -801
rect -1513 -1198 -1475 -801
rect -1347 -1198 -1309 -801
rect -1181 -1198 -1143 -801
rect -1015 -1198 -977 -801
rect -849 -1198 -811 -801
rect -683 -1198 -645 -801
rect -517 -1198 -479 -801
rect -351 -1198 -313 -801
rect -185 -1198 -147 -801
rect -19 -1198 19 -801
rect 147 -1198 185 -801
rect 313 -1198 351 -801
rect 479 -1198 517 -801
rect 645 -1198 683 -801
rect 811 -1198 849 -801
rect 977 -1198 1015 -801
rect 1143 -1198 1181 -801
rect 1309 -1198 1347 -801
rect 1475 -1198 1513 -801
rect 1641 -1198 1679 -801
rect 1807 -1198 1845 -801
rect 1973 -1198 2011 -801
<< metal1 >>
rect -2017 1198 -1967 1210
rect -2017 801 -2011 1198
rect -1973 801 -1967 1198
rect -2017 789 -1967 801
rect -1851 1198 -1801 1210
rect -1851 801 -1845 1198
rect -1807 801 -1801 1198
rect -1851 789 -1801 801
rect -1685 1198 -1635 1210
rect -1685 801 -1679 1198
rect -1641 801 -1635 1198
rect -1685 789 -1635 801
rect -1519 1198 -1469 1210
rect -1519 801 -1513 1198
rect -1475 801 -1469 1198
rect -1519 789 -1469 801
rect -1353 1198 -1303 1210
rect -1353 801 -1347 1198
rect -1309 801 -1303 1198
rect -1353 789 -1303 801
rect -1187 1198 -1137 1210
rect -1187 801 -1181 1198
rect -1143 801 -1137 1198
rect -1187 789 -1137 801
rect -1021 1198 -971 1210
rect -1021 801 -1015 1198
rect -977 801 -971 1198
rect -1021 789 -971 801
rect -855 1198 -805 1210
rect -855 801 -849 1198
rect -811 801 -805 1198
rect -855 789 -805 801
rect -689 1198 -639 1210
rect -689 801 -683 1198
rect -645 801 -639 1198
rect -689 789 -639 801
rect -523 1198 -473 1210
rect -523 801 -517 1198
rect -479 801 -473 1198
rect -523 789 -473 801
rect -357 1198 -307 1210
rect -357 801 -351 1198
rect -313 801 -307 1198
rect -357 789 -307 801
rect -191 1198 -141 1210
rect -191 801 -185 1198
rect -147 801 -141 1198
rect -191 789 -141 801
rect -25 1198 25 1210
rect -25 801 -19 1198
rect 19 801 25 1198
rect -25 789 25 801
rect 141 1198 191 1210
rect 141 801 147 1198
rect 185 801 191 1198
rect 141 789 191 801
rect 307 1198 357 1210
rect 307 801 313 1198
rect 351 801 357 1198
rect 307 789 357 801
rect 473 1198 523 1210
rect 473 801 479 1198
rect 517 801 523 1198
rect 473 789 523 801
rect 639 1198 689 1210
rect 639 801 645 1198
rect 683 801 689 1198
rect 639 789 689 801
rect 805 1198 855 1210
rect 805 801 811 1198
rect 849 801 855 1198
rect 805 789 855 801
rect 971 1198 1021 1210
rect 971 801 977 1198
rect 1015 801 1021 1198
rect 971 789 1021 801
rect 1137 1198 1187 1210
rect 1137 801 1143 1198
rect 1181 801 1187 1198
rect 1137 789 1187 801
rect 1303 1198 1353 1210
rect 1303 801 1309 1198
rect 1347 801 1353 1198
rect 1303 789 1353 801
rect 1469 1198 1519 1210
rect 1469 801 1475 1198
rect 1513 801 1519 1198
rect 1469 789 1519 801
rect 1635 1198 1685 1210
rect 1635 801 1641 1198
rect 1679 801 1685 1198
rect 1635 789 1685 801
rect 1801 1198 1851 1210
rect 1801 801 1807 1198
rect 1845 801 1851 1198
rect 1801 789 1851 801
rect 1967 1198 2017 1210
rect 1967 801 1973 1198
rect 2011 801 2017 1198
rect 1967 789 2017 801
rect -2017 -801 -1967 -789
rect -2017 -1198 -2011 -801
rect -1973 -1198 -1967 -801
rect -2017 -1210 -1967 -1198
rect -1851 -801 -1801 -789
rect -1851 -1198 -1845 -801
rect -1807 -1198 -1801 -801
rect -1851 -1210 -1801 -1198
rect -1685 -801 -1635 -789
rect -1685 -1198 -1679 -801
rect -1641 -1198 -1635 -801
rect -1685 -1210 -1635 -1198
rect -1519 -801 -1469 -789
rect -1519 -1198 -1513 -801
rect -1475 -1198 -1469 -801
rect -1519 -1210 -1469 -1198
rect -1353 -801 -1303 -789
rect -1353 -1198 -1347 -801
rect -1309 -1198 -1303 -801
rect -1353 -1210 -1303 -1198
rect -1187 -801 -1137 -789
rect -1187 -1198 -1181 -801
rect -1143 -1198 -1137 -801
rect -1187 -1210 -1137 -1198
rect -1021 -801 -971 -789
rect -1021 -1198 -1015 -801
rect -977 -1198 -971 -801
rect -1021 -1210 -971 -1198
rect -855 -801 -805 -789
rect -855 -1198 -849 -801
rect -811 -1198 -805 -801
rect -855 -1210 -805 -1198
rect -689 -801 -639 -789
rect -689 -1198 -683 -801
rect -645 -1198 -639 -801
rect -689 -1210 -639 -1198
rect -523 -801 -473 -789
rect -523 -1198 -517 -801
rect -479 -1198 -473 -801
rect -523 -1210 -473 -1198
rect -357 -801 -307 -789
rect -357 -1198 -351 -801
rect -313 -1198 -307 -801
rect -357 -1210 -307 -1198
rect -191 -801 -141 -789
rect -191 -1198 -185 -801
rect -147 -1198 -141 -801
rect -191 -1210 -141 -1198
rect -25 -801 25 -789
rect -25 -1198 -19 -801
rect 19 -1198 25 -801
rect -25 -1210 25 -1198
rect 141 -801 191 -789
rect 141 -1198 147 -801
rect 185 -1198 191 -801
rect 141 -1210 191 -1198
rect 307 -801 357 -789
rect 307 -1198 313 -801
rect 351 -1198 357 -801
rect 307 -1210 357 -1198
rect 473 -801 523 -789
rect 473 -1198 479 -801
rect 517 -1198 523 -801
rect 473 -1210 523 -1198
rect 639 -801 689 -789
rect 639 -1198 645 -801
rect 683 -1198 689 -801
rect 639 -1210 689 -1198
rect 805 -801 855 -789
rect 805 -1198 811 -801
rect 849 -1198 855 -801
rect 805 -1210 855 -1198
rect 971 -801 1021 -789
rect 971 -1198 977 -801
rect 1015 -1198 1021 -801
rect 971 -1210 1021 -1198
rect 1137 -801 1187 -789
rect 1137 -1198 1143 -801
rect 1181 -1198 1187 -801
rect 1137 -1210 1187 -1198
rect 1303 -801 1353 -789
rect 1303 -1198 1309 -801
rect 1347 -1198 1353 -801
rect 1303 -1210 1353 -1198
rect 1469 -801 1519 -789
rect 1469 -1198 1475 -801
rect 1513 -1198 1519 -801
rect 1469 -1210 1519 -1198
rect 1635 -801 1685 -789
rect 1635 -1198 1641 -801
rect 1679 -1198 1685 -801
rect 1635 -1210 1685 -1198
rect 1801 -801 1851 -789
rect 1801 -1198 1807 -801
rect 1845 -1198 1851 -801
rect 1801 -1210 1851 -1198
rect 1967 -801 2017 -789
rect 1967 -1198 1973 -801
rect 2011 -1198 2017 -801
rect 1967 -1210 2017 -1198
<< properties >>
string FIXED_BBOX -2140 -1329 2140 1329
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 8.0 m 1 nx 25 wmin 0.350 lmin 0.50 rho 2000 val 46.789k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
