VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__xtal_osc_16M
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__xtal_osc_16M ;
  ORIGIN 0.000 0.000 ;
  SIZE 54.520 BY 28.480 ;
  PIN in
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.526800 ;
    PORT
      LAYER met1 ;
        RECT 0.000 17.280 1.000 18.280 ;
    END
  END in
  PIN out
    PORT
      LAYER met1 ;
        RECT 0.000 8.590 1.000 9.590 ;
    END
  END out
  PIN avdd
    ANTENNADIFFAREA 98.890800 ;
    PORT
      LAYER met2 ;
        RECT 0.000 20.135 0.625 28.275 ;
    END
  END avdd
  PIN avss
    ANTENNADIFFAREA 87.223801 ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.125 4.565 8.250 ;
    END
  END avss
  PIN dvdd
    ANTENNADIFFAREA 4.959600 ;
    PORT
      LAYER met2 ;
        RECT 53.615 14.290 54.520 18.150 ;
    END
  END dvdd
  PIN dvss
    ANTENNADIFFAREA 21.305099 ;
    PORT
      LAYER met1 ;
        RECT 53.395 0.460 54.520 5.280 ;
    END
  END dvss
  PIN ena
    ANTENNAGATEAREA 0.510000 ;
    PORT
      LAYER met1 ;
        RECT 52.670 7.390 54.520 8.390 ;
    END
  END ena
  PIN dout
    ANTENNADIFFAREA 0.435000 ;
    PORT
      LAYER met1 ;
        RECT 53.520 12.640 54.520 13.640 ;
    END
  END dout
  PIN stdby
    ANTENNAGATEAREA 0.510000 ;
    PORT
      LAYER met1 ;
        RECT 52.670 20.070 54.520 21.070 ;
    END
  END stdby
  OBS
      LAYER nwell ;
        RECT 0.000 26.870 47.350 28.480 ;
        RECT 0.000 1.590 1.610 26.870 ;
        RECT 0.000 0.000 47.350 1.590 ;
      LAYER li1 ;
        RECT 0.465 0.420 54.510 28.015 ;
      LAYER met1 ;
        RECT 0.530 21.350 54.520 28.045 ;
        RECT 0.530 19.790 52.390 21.350 ;
        RECT 0.530 18.560 54.520 19.790 ;
        RECT 1.280 17.000 54.520 18.560 ;
        RECT 0.530 13.920 54.520 17.000 ;
        RECT 0.530 12.360 53.240 13.920 ;
        RECT 0.530 9.870 54.520 12.360 ;
        RECT 1.280 8.670 54.520 9.870 ;
        RECT 1.280 8.310 52.390 8.670 ;
        RECT 0.530 7.110 52.390 8.310 ;
        RECT 0.530 5.560 54.520 7.110 ;
        RECT 0.530 0.420 53.115 5.560 ;
      LAYER met2 ;
        RECT 0.905 19.855 53.685 28.285 ;
        RECT 0.625 18.430 53.685 19.855 ;
        RECT 0.625 14.010 53.335 18.430 ;
        RECT 0.625 8.530 53.685 14.010 ;
        RECT 4.845 0.125 53.685 8.530 ;
  END
END sky130_ef_ip__xtal_osc_16M
END LIBRARY

