magic
tech sky130A
magscale 1 2
timestamp 1698886478
<< pwell >>
rect -948 -1382 948 1382
<< psubdiff >>
rect -912 1312 -816 1346
rect 816 1312 912 1346
rect -912 1250 -878 1312
rect 878 1250 912 1312
rect -912 -1312 -878 -1250
rect 878 -1312 912 -1250
rect -912 -1346 -816 -1312
rect 816 -1346 912 -1312
<< psubdiffcont >>
rect -816 1312 816 1346
rect -912 -1250 -878 1250
rect 878 -1250 912 1250
rect -816 -1346 816 -1312
<< xpolycontact >>
rect -782 784 -712 1216
rect -782 -1216 -712 -784
rect -616 784 -546 1216
rect -616 -1216 -546 -784
rect -450 784 -380 1216
rect -450 -1216 -380 -784
rect -284 784 -214 1216
rect -284 -1216 -214 -784
rect -118 784 -48 1216
rect -118 -1216 -48 -784
rect 48 784 118 1216
rect 48 -1216 118 -784
rect 214 784 284 1216
rect 214 -1216 284 -784
rect 380 784 450 1216
rect 380 -1216 450 -784
rect 546 784 616 1216
rect 546 -1216 616 -784
rect 712 784 782 1216
rect 712 -1216 782 -784
<< xpolyres >>
rect -782 -784 -712 784
rect -616 -784 -546 784
rect -450 -784 -380 784
rect -284 -784 -214 784
rect -118 -784 -48 784
rect 48 -784 118 784
rect 214 -784 284 784
rect 380 -784 450 784
rect 546 -784 616 784
rect 712 -784 782 784
<< locali >>
rect -912 1312 -816 1346
rect 816 1312 912 1346
rect -912 1250 -878 1312
rect 878 1250 912 1312
rect -912 -1312 -878 -1250
rect 878 -1312 912 -1250
rect -912 -1346 -816 -1312
rect 816 -1346 912 -1312
<< viali >>
rect -766 801 -728 1198
rect -600 801 -562 1198
rect -434 801 -396 1198
rect -268 801 -230 1198
rect -102 801 -64 1198
rect 64 801 102 1198
rect 230 801 268 1198
rect 396 801 434 1198
rect 562 801 600 1198
rect 728 801 766 1198
rect -766 -1198 -728 -801
rect -600 -1198 -562 -801
rect -434 -1198 -396 -801
rect -268 -1198 -230 -801
rect -102 -1198 -64 -801
rect 64 -1198 102 -801
rect 230 -1198 268 -801
rect 396 -1198 434 -801
rect 562 -1198 600 -801
rect 728 -1198 766 -801
<< metal1 >>
rect -772 1198 -722 1210
rect -772 801 -766 1198
rect -728 801 -722 1198
rect -772 789 -722 801
rect -606 1198 -556 1210
rect -606 801 -600 1198
rect -562 801 -556 1198
rect -606 789 -556 801
rect -440 1198 -390 1210
rect -440 801 -434 1198
rect -396 801 -390 1198
rect -440 789 -390 801
rect -274 1198 -224 1210
rect -274 801 -268 1198
rect -230 801 -224 1198
rect -274 789 -224 801
rect -108 1198 -58 1210
rect -108 801 -102 1198
rect -64 801 -58 1198
rect -108 789 -58 801
rect 58 1198 108 1210
rect 58 801 64 1198
rect 102 801 108 1198
rect 58 789 108 801
rect 224 1198 274 1210
rect 224 801 230 1198
rect 268 801 274 1198
rect 224 789 274 801
rect 390 1198 440 1210
rect 390 801 396 1198
rect 434 801 440 1198
rect 390 789 440 801
rect 556 1198 606 1210
rect 556 801 562 1198
rect 600 801 606 1198
rect 556 789 606 801
rect 722 1198 772 1210
rect 722 801 728 1198
rect 766 801 772 1198
rect 722 789 772 801
rect -772 -801 -722 -789
rect -772 -1198 -766 -801
rect -728 -1198 -722 -801
rect -772 -1210 -722 -1198
rect -606 -801 -556 -789
rect -606 -1198 -600 -801
rect -562 -1198 -556 -801
rect -606 -1210 -556 -1198
rect -440 -801 -390 -789
rect -440 -1198 -434 -801
rect -396 -1198 -390 -801
rect -440 -1210 -390 -1198
rect -274 -801 -224 -789
rect -274 -1198 -268 -801
rect -230 -1198 -224 -801
rect -274 -1210 -224 -1198
rect -108 -801 -58 -789
rect -108 -1198 -102 -801
rect -64 -1198 -58 -801
rect -108 -1210 -58 -1198
rect 58 -801 108 -789
rect 58 -1198 64 -801
rect 102 -1198 108 -801
rect 58 -1210 108 -1198
rect 224 -801 274 -789
rect 224 -1198 230 -801
rect 268 -1198 274 -801
rect 224 -1210 274 -1198
rect 390 -801 440 -789
rect 390 -1198 396 -801
rect 434 -1198 440 -801
rect 390 -1210 440 -1198
rect 556 -801 606 -789
rect 556 -1198 562 -801
rect 600 -1198 606 -801
rect 556 -1210 606 -1198
rect 722 -801 772 -789
rect 722 -1198 728 -801
rect 766 -1198 772 -801
rect 722 -1210 772 -1198
<< properties >>
string FIXED_BBOX -895 -1329 895 1329
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 8.0 m 1 nx 10 wmin 0.350 lmin 0.50 rho 2000 val 46.789k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
