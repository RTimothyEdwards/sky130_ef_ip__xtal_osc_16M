magic
tech sky130A
magscale 1 2
timestamp 1699037441
<< dnwell >>
rect 2576 -2328 11814 3140
<< nwell >>
rect 2460 2934 11930 3256
rect 2460 -2122 2782 2934
rect 11608 -2122 11930 2934
rect 2460 -2440 11930 -2122
<< psubdiff >>
rect 12438 3146 13362 3151
rect 12438 3108 12508 3146
rect 13295 3108 13362 3146
rect 12438 3101 13362 3108
rect 12438 3056 12488 3101
rect 12438 -2243 12447 3056
rect 12481 -2243 12488 3056
rect 12438 -2306 12488 -2243
rect 13312 3056 13362 3101
rect 13312 -2243 13321 3056
rect 13355 -2243 13362 3056
rect 13312 -2306 13362 -2243
rect 12438 -2312 13362 -2306
rect 12438 -2350 12515 -2312
rect 13302 -2350 13362 -2312
rect 12438 -2356 13362 -2350
<< mvnsubdiff >>
rect 2533 3163 11857 3183
rect 2533 3129 2613 3163
rect 11777 3129 11857 3163
rect 2533 3109 11857 3129
rect 2533 3103 2607 3109
rect 2533 -2291 2553 3103
rect 2587 -2291 2607 3103
rect 2533 -2297 2607 -2291
rect 11783 3103 11857 3109
rect 11783 -2291 11803 3103
rect 11837 -2291 11857 3103
rect 11783 -2297 11857 -2291
rect 2533 -2317 11857 -2297
rect 2533 -2351 2613 -2317
rect 11777 -2351 11857 -2317
rect 2533 -2371 11857 -2351
<< psubdiffcont >>
rect 12508 3108 13295 3146
rect 12447 -2243 12481 3056
rect 13321 -2243 13355 3056
rect 12515 -2350 13302 -2312
<< mvnsubdiffcont >>
rect 2613 3129 11777 3163
rect 2553 -2291 2587 3103
rect 11803 -2291 11837 3103
rect 2613 -2351 11777 -2317
<< locali >>
rect 2553 3129 2613 3163
rect 11777 3140 12035 3163
rect 11777 3129 11860 3140
rect 2553 3114 2693 3129
rect 2553 3103 2585 3114
rect 2668 1605 2693 3114
rect 11803 3103 11860 3129
rect 2830 2982 10050 3000
rect 2830 2926 2870 2982
rect 4698 2976 10050 2982
rect 4698 2926 5034 2976
rect 9959 2926 10050 2976
rect 2830 2862 10050 2926
rect 2830 2855 7100 2862
rect 2830 2852 4733 2855
rect 2587 861 2693 1605
rect 2663 131 2693 861
rect 4644 232 4733 2852
rect 4596 228 4733 232
rect 2587 -863 2693 131
rect 2832 126 4733 228
rect 4937 2852 7100 2855
rect 7545 2852 10050 2862
rect 4937 232 5028 2852
rect 9299 1817 9438 2852
rect 9299 240 9334 1817
rect 9401 240 9438 1817
rect 4937 228 5057 232
rect 9299 228 9438 240
rect 9524 2244 9663 2852
rect 9524 247 9557 2244
rect 9624 247 9663 2244
rect 9524 228 9663 247
rect 4937 224 7100 228
rect 7545 224 9667 228
rect 4937 126 9667 224
rect 2832 86 9667 126
rect 2832 17 3549 86
rect 2553 -2313 2581 -2291
rect 2662 -2313 2693 -863
rect 3299 -52 3549 17
rect 3299 -2018 3373 -52
rect 3483 -171 3549 -52
rect 4009 9 8864 14
rect 4009 4 6477 9
rect 4009 -126 5294 4
rect 5934 -121 6477 4
rect 7117 7 8864 9
rect 7117 -121 7624 7
rect 5934 -126 7624 -121
rect 4009 -129 7624 -126
rect 8023 -129 8864 7
rect 4009 -140 8864 -129
rect 8958 -1 9667 86
rect 3483 -284 3899 -171
rect 3483 -533 3549 -284
rect 3814 -533 3899 -284
rect 3483 -909 3899 -533
rect 4009 -590 4130 -140
rect 4009 -592 4418 -590
rect 4009 -740 4100 -592
rect 4240 -740 4418 -592
rect 4860 -592 8870 -590
rect 4860 -740 5164 -592
rect 4009 -741 5164 -740
rect 6078 -594 8870 -592
rect 6078 -741 6344 -594
rect 6699 -741 6965 -594
rect 7320 -741 8870 -594
rect 4009 -744 8870 -741
rect 3483 -910 3818 -909
rect 3483 -2018 3549 -910
rect 3299 -2054 3549 -2018
rect 3300 -2060 3549 -2054
rect 4545 -976 8406 -816
rect 4545 -1406 4643 -976
rect 4545 -1421 8408 -1406
rect 4545 -1422 7466 -1421
rect 4545 -1560 4621 -1422
rect 4768 -1560 5199 -1422
rect 5346 -1424 6835 -1422
rect 5346 -1560 5760 -1424
rect 4545 -1562 5760 -1560
rect 5907 -1560 6835 -1424
rect 6982 -1559 7466 -1422
rect 8289 -1559 8408 -1421
rect 6982 -1560 8408 -1559
rect 5907 -1562 8408 -1560
rect 4545 -1566 8408 -1562
rect 4545 -2004 4643 -1566
rect 4545 -2023 8400 -2004
rect 4545 -2144 4622 -2023
rect 8372 -2144 8400 -2023
rect 4545 -2164 8400 -2144
rect 8958 -2027 9058 -1
rect 9510 -20 9667 -1
rect 9496 -105 9669 -20
rect 9496 -521 9501 -105
rect 9603 -177 9669 -105
rect 9945 -177 10046 2852
rect 9603 -323 10046 -177
rect 9603 -521 9669 -323
rect 9496 -1179 9669 -521
rect 9495 -1192 9768 -1179
rect 9495 -1565 9505 -1192
rect 9756 -1565 9768 -1192
rect 9495 -1577 9768 -1565
rect 9496 -1874 9669 -1577
rect 9496 -1887 9975 -1874
rect 9496 -2027 9509 -1887
rect 8958 -2188 9509 -2027
rect 9496 -2222 9509 -2188
rect 9963 -2222 9975 -1887
rect 9496 -2236 9975 -2222
rect 2553 -2317 2693 -2313
rect 11837 -2291 11860 3103
rect 11803 -2317 11860 -2291
rect 2553 -2351 2613 -2317
rect 11777 -2323 11860 -2317
rect 12024 -2323 12035 3140
rect 11777 -2351 12035 -2323
rect 12261 3146 13362 3151
rect 12261 3132 12508 3146
rect 12261 -2315 12290 3132
rect 12422 3108 12508 3132
rect 13295 3108 13362 3146
rect 12422 3056 13362 3108
rect 12422 -2243 12447 3056
rect 12481 3037 13321 3056
rect 12481 2859 12580 3037
rect 13247 2859 13321 3037
rect 12481 2197 13321 2859
rect 12481 1731 12753 2197
rect 12481 36 12488 1731
rect 12655 870 13250 886
rect 12655 808 12958 870
rect 13116 808 13250 870
rect 12655 785 13250 808
rect 12655 467 12790 785
rect 13312 346 13321 2197
rect 13016 324 13321 346
rect 12481 28 12667 36
rect 13021 28 13321 324
rect 12481 12 13321 28
rect 12481 -37 12515 12
rect 12873 -37 13321 12
rect 12481 -78 13321 -37
rect 12481 -918 12488 -78
rect 12481 -1410 12768 -918
rect 13312 -1410 13321 -78
rect 12481 -2076 13321 -1410
rect 12481 -2243 12571 -2076
rect 12422 -2254 12571 -2243
rect 13139 -2243 13321 -2076
rect 13355 -2243 13362 3056
rect 13139 -2254 13362 -2243
rect 12422 -2312 13362 -2254
rect 12422 -2315 12515 -2312
rect 12261 -2350 12515 -2315
rect 13302 -2350 13362 -2312
rect 12261 -2356 13362 -2350
<< viali >>
rect 2585 3103 2668 3114
rect 2585 1605 2587 3103
rect 2587 1605 2668 3103
rect 2870 2926 4698 2982
rect 5034 2926 9959 2976
rect 2581 131 2587 861
rect 2587 131 2663 861
rect 4733 126 4937 2855
rect 9334 240 9401 1817
rect 9557 247 9624 2244
rect 2581 -2291 2587 -863
rect 2587 -2291 2662 -863
rect 2581 -2313 2662 -2291
rect 3373 -2018 3483 -52
rect 5294 -126 5934 4
rect 6477 -121 7117 9
rect 7624 -129 8023 7
rect 4100 -740 4240 -592
rect 4418 -740 4860 -590
rect 5164 -741 6078 -592
rect 6344 -741 6699 -594
rect 6965 -741 7320 -594
rect 4621 -1560 4768 -1422
rect 5199 -1560 5346 -1422
rect 5760 -1562 5907 -1424
rect 6835 -1560 6982 -1422
rect 7466 -1559 8289 -1421
rect 4622 -2144 8372 -2023
rect 9501 -521 9603 -105
rect 9505 -1565 9756 -1192
rect 9509 -2222 9963 -1887
rect 11860 -2323 12024 3140
rect 12290 -2315 12422 3132
rect 12580 2859 13247 3037
rect 12958 808 13116 870
rect 12515 -37 12873 12
rect 12571 -2254 13139 -2076
<< metal1 >>
rect 2579 3114 2674 3126
rect 2575 1605 2585 3114
rect 2668 1605 2678 3114
rect 2801 2982 11608 2999
rect 2801 2926 2870 2982
rect 4698 2976 11608 2982
rect 4698 2926 5034 2976
rect 9959 2926 11608 2976
rect 2801 2855 11608 2926
rect 2801 2854 4733 2855
rect 2964 2328 3200 2760
rect 3296 2328 3532 2760
rect 3628 2328 3864 2760
rect 3960 2328 4196 2760
rect 4292 2328 4528 2760
rect 2579 1593 2674 1605
rect 2460 1128 2660 1216
rect 2460 1093 2774 1128
rect 2460 1016 2660 1093
rect 2569 861 2680 882
rect 2569 131 2581 861
rect 2663 131 2680 861
rect 2569 114 2680 131
rect 2739 67 2774 1093
rect 2838 746 3034 760
rect 2838 345 2852 746
rect 3015 345 3034 746
rect 2838 328 3034 345
rect 3130 328 3366 760
rect 3462 328 3698 760
rect 3794 328 4030 760
rect 4126 328 4362 760
rect 4472 384 4509 402
rect 4472 329 4520 384
rect 3096 139 3106 204
rect 3307 139 3317 204
rect 2721 2 2731 67
rect 2932 2 2942 67
rect 3136 -121 3179 139
rect 4472 122 4509 329
rect 3947 85 4509 122
rect 4694 126 4733 2854
rect 4937 2854 11608 2855
rect 4937 126 4983 2854
rect 5134 2327 5370 2759
rect 5466 2327 5702 2759
rect 5798 2327 6034 2759
rect 6130 2327 6366 2759
rect 6462 2327 6698 2759
rect 6794 2327 7030 2759
rect 7126 2327 7362 2759
rect 7458 2327 7694 2759
rect 7790 2327 8026 2759
rect 8122 2327 8358 2759
rect 8454 2327 8690 2759
rect 8786 2327 9022 2759
rect 9118 2393 9188 2759
rect 9428 2753 9837 2759
rect 9118 2349 9393 2393
rect 9118 2326 9188 2349
rect 9349 2104 9393 2349
rect 9428 2330 9452 2753
rect 9624 2330 9837 2753
rect 9428 2326 9837 2330
rect 9551 2255 9630 2256
rect 9542 2244 9638 2255
rect 9329 1898 9339 2104
rect 9397 1898 9407 2104
rect 9320 1817 9416 1832
rect 5134 695 5182 745
rect 5141 327 5195 403
rect 5300 327 5536 759
rect 5632 327 5868 759
rect 5964 327 6200 759
rect 6296 327 6532 759
rect 6628 327 6864 759
rect 6960 327 7196 759
rect 7292 327 7528 759
rect 7624 327 7860 759
rect 7956 327 8192 759
rect 8288 327 8524 759
rect 8620 327 8856 759
rect 8952 327 9188 759
rect 4694 105 4983 126
rect 3563 4 3573 69
rect 3774 4 3784 69
rect 3358 -52 3493 -38
rect 2460 -579 2660 -522
rect 2460 -640 2874 -579
rect 2460 -722 2660 -640
rect 2566 -863 2678 -846
rect 2566 -2313 2581 -863
rect 2662 -2313 2678 -863
rect 2813 -1507 2874 -640
rect 2813 -1568 3188 -1507
rect 3358 -2018 3373 -52
rect 3483 -2018 3493 -52
rect 3657 -667 3704 4
rect 3657 -714 3841 -667
rect 3794 -1197 3841 -714
rect 3947 -1167 3984 85
rect 5147 56 5185 327
rect 9118 326 9188 327
rect 9320 240 9334 1817
rect 9401 240 9416 1817
rect 7183 230 7629 231
rect 5278 228 6454 229
rect 7183 228 8031 230
rect 5278 221 8031 228
rect 9320 224 9416 240
rect 9542 247 9557 2244
rect 9624 247 9638 2244
rect 11719 2202 11744 3169
rect 12055 2202 12077 3169
rect 9542 227 9638 247
rect 10040 1342 10162 1378
rect 5278 214 7451 221
rect 5278 115 6445 214
rect 4987 -9 4997 56
rect 5198 -9 5208 56
rect 5278 4 5947 115
rect 5278 -126 5294 4
rect 5934 -126 5947 4
rect 5994 3 6004 68
rect 6205 3 6215 68
rect 5278 -127 5947 -126
rect 5282 -132 5946 -127
rect 4163 -580 4244 -323
rect 4094 -592 4246 -580
rect 4090 -740 4100 -592
rect 4240 -740 4250 -592
rect 4094 -752 4246 -740
rect 4307 -1049 4343 -238
rect 4404 -272 5605 -234
rect 4404 -412 4442 -272
rect 4781 -584 4862 -323
rect 4926 -479 4958 -272
rect 4406 -590 4872 -584
rect 4406 -740 4418 -590
rect 4860 -740 4872 -590
rect 4406 -746 4872 -740
rect 5032 -909 5078 -272
rect 5397 -586 5478 -325
rect 5537 -480 5569 -272
rect 5641 -385 6095 -349
rect 5152 -592 6090 -586
rect 5152 -741 5164 -592
rect 6078 -741 6090 -592
rect 5152 -747 6090 -741
rect 5032 -955 5526 -909
rect 6163 -933 6198 3
rect 6424 -39 6445 115
rect 7229 -31 7451 214
rect 8011 13 8031 221
rect 8244 112 8254 177
rect 8455 112 8465 177
rect 8515 123 9789 157
rect 8011 7 8035 13
rect 7229 -39 7624 -31
rect 6424 -121 6477 -39
rect 7117 -74 7624 -39
rect 7117 -121 7250 -74
rect 6424 -127 7250 -121
rect 6424 -321 6700 -127
rect 6257 -871 6299 -323
rect 6424 -588 6701 -321
rect 6332 -594 6711 -588
rect 6332 -741 6344 -594
rect 6699 -741 6711 -594
rect 6332 -747 6711 -741
rect 6776 -871 6813 -248
rect 6986 -319 7250 -127
rect 7335 -191 7345 -126
rect 7546 -191 7556 -126
rect 7604 -129 7624 -74
rect 8023 -129 8035 7
rect 8165 -7 8175 22
rect 7604 -135 8035 -129
rect 8114 -43 8175 -7
rect 8376 -43 8386 22
rect 7604 -136 8031 -135
rect 6869 -777 6906 -323
rect 6986 -588 7326 -319
rect 6953 -594 7332 -588
rect 6953 -741 6965 -594
rect 7320 -741 7332 -594
rect 6953 -747 7332 -741
rect 6869 -782 7187 -777
rect 7395 -782 7431 -253
rect 7495 -656 7535 -191
rect 7713 -412 7723 -319
rect 7965 -412 7975 -319
rect 7495 -696 7745 -656
rect 6869 -814 7636 -782
rect 7150 -818 7636 -814
rect 6257 -908 7084 -871
rect 5990 -954 6000 -933
rect 4237 -1114 4247 -1049
rect 4448 -1114 4458 -1049
rect 5002 -1072 5012 -1055
rect 4817 -1108 5012 -1072
rect 3947 -1204 4767 -1167
rect 4820 -1290 4858 -1108
rect 5002 -1120 5012 -1108
rect 5213 -1072 5223 -1055
rect 5213 -1108 5410 -1072
rect 5213 -1120 5223 -1108
rect 4609 -1422 4780 -1416
rect 4609 -1560 4621 -1422
rect 4768 -1560 4780 -1422
rect 4609 -1566 4780 -1560
rect 4696 -1832 4756 -1566
rect 4818 -1898 4854 -1698
rect 4924 -1898 4968 -1140
rect 5268 -1342 5312 -1142
rect 5372 -1296 5410 -1108
rect 5480 -1230 5526 -955
rect 5934 -998 6000 -954
rect 6201 -998 6211 -933
rect 5822 -1340 5866 -1146
rect 5934 -1302 5969 -998
rect 6257 -1152 6299 -908
rect 6031 -1194 6300 -1152
rect 6031 -1235 6073 -1194
rect 5268 -1386 5528 -1342
rect 5822 -1384 6082 -1340
rect 5187 -1422 5358 -1416
rect 5187 -1560 5199 -1422
rect 5346 -1560 5358 -1422
rect 5187 -1566 5358 -1560
rect 5244 -1830 5304 -1566
rect 5378 -1898 5414 -1692
rect 5484 -1832 5528 -1386
rect 5748 -1424 5919 -1418
rect 5748 -1562 5760 -1424
rect 5907 -1562 5919 -1424
rect 5748 -1568 5919 -1562
rect 5808 -1832 5868 -1568
rect 5934 -1894 5970 -1686
rect 6038 -1834 6082 -1384
rect 6907 -1416 6984 -1146
rect 7047 -1274 7084 -908
rect 7150 -1235 7187 -818
rect 7266 -1003 7276 -938
rect 7477 -1003 7487 -938
rect 6823 -1422 6994 -1416
rect 6823 -1560 6835 -1422
rect 6982 -1560 6994 -1422
rect 7042 -1470 7085 -1274
rect 7042 -1513 7194 -1470
rect 6823 -1566 6994 -1560
rect 6907 -1570 6984 -1566
rect 6492 -1656 6526 -1654
rect 6680 -1656 6690 -1643
rect 6484 -1694 6690 -1656
rect 6213 -1811 6435 -1771
rect 6213 -1898 6253 -1811
rect 6492 -1893 6526 -1694
rect 6680 -1708 6690 -1694
rect 6891 -1656 6901 -1643
rect 6891 -1694 7108 -1656
rect 6891 -1708 6901 -1694
rect 4796 -1938 6253 -1898
rect 6593 -2005 6665 -1742
rect 6900 -2005 6983 -1750
rect 7045 -1896 7079 -1694
rect 7151 -1837 7194 -1513
rect 7335 -1772 7375 -1003
rect 7466 -1415 7543 -1142
rect 7600 -1277 7636 -818
rect 7705 -1233 7745 -696
rect 8005 -785 8037 -258
rect 8114 -691 8150 -43
rect 8414 -381 8446 112
rect 8364 -413 8446 -381
rect 8515 -411 8549 123
rect 8616 17 9714 53
rect 8114 -727 8295 -691
rect 8005 -817 8190 -785
rect 8158 -1064 8190 -817
rect 7860 -1100 8191 -1064
rect 7860 -1277 7896 -1100
rect 7600 -1313 7896 -1277
rect 8010 -1415 8087 -1141
rect 8158 -1298 8190 -1100
rect 8259 -1236 8295 -727
rect 7454 -1421 8301 -1415
rect 7454 -1559 7466 -1421
rect 8289 -1559 8301 -1421
rect 7454 -1565 8301 -1559
rect 7466 -1566 7543 -1565
rect 7582 -1646 8224 -1642
rect 8364 -1646 8396 -413
rect 8616 -464 8652 17
rect 9495 -98 9609 -93
rect 9329 -105 9610 -98
rect 8737 -336 9179 -323
rect 8716 -388 9186 -336
rect 8737 -391 9179 -388
rect 8471 -560 8511 -551
rect 8464 -625 8474 -560
rect 8675 -625 8685 -560
rect 7582 -1678 8396 -1646
rect 7582 -1686 8224 -1678
rect 7335 -1812 7551 -1772
rect 7596 -1907 7634 -1688
rect 7707 -1937 7790 -1749
rect 8012 -1937 8095 -1751
rect 8157 -1898 8195 -1686
rect 8471 -1769 8511 -625
rect 8737 -712 8805 -391
rect 9329 -521 9501 -105
rect 9603 -521 9610 -105
rect 9678 -138 9714 17
rect 10040 -138 10076 1342
rect 10104 1123 10114 1188
rect 10315 1123 10325 1188
rect 11719 637 11860 2202
rect 11597 -40 11860 637
rect 9678 -174 10076 -138
rect 10106 -372 10116 -307
rect 10317 -372 10327 -307
rect 9329 -531 9610 -521
rect 9495 -533 9609 -531
rect 10106 -599 10116 -534
rect 10317 -599 10327 -534
rect 8244 -1809 8511 -1769
rect 8554 -780 8805 -712
rect 7707 -1938 8095 -1937
rect 8554 -1938 8622 -780
rect 9495 -1192 9768 -1179
rect 9163 -1931 9399 -1499
rect 9495 -1565 9505 -1192
rect 9756 -1565 9768 -1192
rect 9495 -1577 9768 -1565
rect 9496 -1886 11684 -1874
rect 9496 -1887 10357 -1886
rect 7707 -1976 8622 -1938
rect 7707 -2005 7790 -2004
rect 8012 -2005 8095 -2004
rect 3358 -2032 3493 -2018
rect 4598 -2023 8401 -2005
rect 4598 -2144 4622 -2023
rect 8372 -2144 8401 -2023
rect 4598 -2164 8401 -2144
rect 9496 -2222 9509 -1887
rect 9963 -2222 10357 -1887
rect 9496 -2224 10357 -2222
rect 11571 -2224 11684 -1886
rect 9496 -2236 11684 -2224
rect 2566 -2331 2678 -2313
rect 11719 -2323 11860 -40
rect 12024 -2323 12077 2202
rect 11719 -2356 12077 -2323
rect 12240 3132 13362 3156
rect 12240 -2315 12290 3132
rect 12422 3037 13362 3132
rect 12422 2859 12580 3037
rect 13247 2859 13362 3037
rect 12422 2196 13362 2859
rect 12422 101 12545 2196
rect 13164 1574 13364 1774
rect 12712 1183 13386 1190
rect 12712 999 12724 1183
rect 13183 999 13386 1183
rect 12712 990 13386 999
rect 12939 870 13142 990
rect 12939 808 12958 870
rect 13116 808 13142 870
rect 12939 694 13142 808
rect 12846 511 12885 675
rect 12770 472 12885 511
rect 12770 427 12809 472
rect 12599 362 12609 427
rect 12810 362 12820 427
rect 12970 413 13014 615
rect 12903 369 13014 413
rect 12770 159 12809 362
rect 12903 268 12947 369
rect 13164 268 13364 288
rect 12903 201 13364 268
rect 12903 200 12947 201
rect 12841 104 12957 122
rect 12840 101 12957 104
rect 12422 12 12959 101
rect 13164 88 13364 201
rect 12422 -37 12515 12
rect 12873 -37 12959 12
rect 12422 -83 12959 -37
rect 12422 -1384 12545 -83
rect 12715 -195 13197 -179
rect 12715 -362 12733 -195
rect 13181 -362 13197 -195
rect 12715 -377 13197 -362
rect 13164 -962 13364 -762
rect 12422 -2076 13364 -1384
rect 12422 -2254 12571 -2076
rect 13139 -2254 13364 -2076
rect 12422 -2315 13364 -2254
rect 12240 -2348 13364 -2315
rect 12240 -2349 12545 -2348
<< via1 >>
rect 2585 1605 2668 3114
rect 2852 345 3015 746
rect 3106 139 3307 204
rect 2731 2 2932 67
rect 9452 2330 9624 2753
rect 9339 1898 9397 2104
rect 3573 4 3774 69
rect 3373 -2018 3481 -805
rect 11744 3140 12055 3169
rect 11744 2202 11860 3140
rect 11860 2202 12024 3140
rect 12024 2202 12055 3140
rect 4997 -9 5198 56
rect 6004 3 6205 68
rect 4100 -740 4240 -592
rect 4418 -740 4860 -590
rect 5164 -741 6078 -592
rect 6445 9 7229 214
rect 6445 -39 6477 9
rect 6477 -39 7117 9
rect 7117 -39 7229 9
rect 7451 7 8011 221
rect 8254 112 8455 177
rect 7451 -31 7624 7
rect 7624 -31 8011 7
rect 6344 -741 6699 -594
rect 7345 -191 7546 -126
rect 8175 -43 8376 22
rect 6965 -741 7320 -594
rect 7723 -412 7965 -319
rect 4247 -1114 4448 -1049
rect 5012 -1120 5213 -1055
rect 4621 -1560 4768 -1422
rect 6000 -998 6201 -933
rect 5199 -1560 5346 -1422
rect 5760 -1562 5907 -1424
rect 7276 -1003 7477 -938
rect 6835 -1560 6982 -1422
rect 6690 -1708 6891 -1643
rect 7466 -1559 8289 -1421
rect 8474 -625 8675 -560
rect 10114 1123 10315 1188
rect 10116 -372 10317 -307
rect 10116 -599 10317 -534
rect 9505 -1565 9756 -1192
rect 4622 -2144 8372 -2023
rect 9509 -2222 9963 -1887
rect 10357 -2224 11571 -1886
rect 12724 999 13183 1183
rect 12609 362 12810 427
rect 12733 -362 13181 -195
<< metal2 >>
rect 9929 3215 12075 3217
rect 2460 3169 12075 3215
rect 2460 3114 11744 3169
rect 2460 1605 2585 3114
rect 2668 2753 11744 3114
rect 2668 2330 9452 2753
rect 9624 2330 11744 2753
rect 2668 2202 11744 2330
rect 12055 2202 12075 3169
rect 2668 2177 12075 2202
rect 2668 1605 9141 2177
rect 9339 2104 9397 2114
rect 9339 1888 9397 1898
rect 2460 1587 9141 1605
rect 2802 746 3056 1587
rect 2802 345 2852 746
rect 3015 345 3056 746
rect 2802 294 3056 345
rect 6426 1213 7256 1587
rect 7420 1213 8033 1587
rect 6426 214 7254 1213
rect 3106 204 3307 214
rect 3307 151 6316 191
rect 3106 129 3307 139
rect 2731 67 2932 77
rect 3573 69 3774 79
rect 2932 17 3573 52
rect 2731 -8 2932 2
rect 6004 68 6205 78
rect 4997 56 5198 66
rect 3774 17 4997 52
rect 3573 -6 3774 4
rect 5198 17 6004 52
rect 6004 -7 6205 3
rect 4997 -19 5198 -9
rect 6276 -139 6316 151
rect 6426 -39 6445 214
rect 7229 -39 7254 214
rect 6426 -56 7254 -39
rect 7422 221 8033 1213
rect 9346 295 9386 1888
rect 10114 1188 10315 1198
rect 7422 -31 7451 221
rect 8011 -31 8033 221
rect 7422 -50 8033 -31
rect 8094 255 9386 295
rect 9854 1125 10114 1175
rect 7345 -126 7546 -116
rect 6276 -179 7345 -139
rect 8094 -139 8134 255
rect 8254 187 8299 188
rect 8254 184 8455 187
rect 9854 184 9904 1125
rect 12712 1183 13386 1190
rect 10315 1125 10378 1175
rect 10114 1113 10315 1123
rect 12712 999 12724 1183
rect 13183 999 13386 1183
rect 12712 990 13386 999
rect 12609 427 12810 437
rect 8254 177 9904 184
rect 8455 134 9904 177
rect 9957 373 12609 417
rect 8254 102 8455 112
rect 9957 52 10001 373
rect 12609 352 12810 362
rect 12888 418 13386 990
rect 8175 22 8376 32
rect 8672 12 10001 52
rect 8376 8 10001 12
rect 8376 -32 8716 8
rect 8175 -53 8376 -43
rect 12888 -54 13196 418
rect 7546 -179 8520 -139
rect 7345 -201 7546 -191
rect 7723 -319 7969 -309
rect 7965 -412 7969 -319
rect 3963 -590 7359 -468
rect 3963 -592 4418 -590
rect 3963 -740 4100 -592
rect 4240 -740 4418 -592
rect 4860 -592 7359 -590
rect 4860 -740 5164 -592
rect 3963 -741 5164 -740
rect 6078 -594 7359 -592
rect 6078 -741 6344 -594
rect 6699 -741 6965 -594
rect 7320 -741 7359 -594
rect 2460 -805 3743 -790
rect 2460 -2018 3373 -805
rect 3481 -1180 3743 -805
rect 3963 -839 7359 -741
rect 7723 -699 7969 -412
rect 8480 -550 8520 -179
rect 8790 -179 13196 -54
rect 8790 -195 13197 -179
rect 8790 -209 12733 -195
rect 8474 -560 8675 -550
rect 8474 -635 8675 -625
rect 8790 -699 8986 -209
rect 10116 -307 10317 -297
rect 7723 -862 8986 -699
rect 9695 -363 10116 -313
rect 6000 -933 6201 -923
rect 7276 -938 7477 -928
rect 6201 -989 7276 -954
rect 6000 -1008 6201 -998
rect 7276 -1013 7477 -1003
rect 4247 -1049 4448 -1039
rect 5012 -1055 5213 -1045
rect 4448 -1109 5012 -1059
rect 4247 -1124 4448 -1114
rect 9695 -1059 9745 -363
rect 10317 -363 10369 -313
rect 12715 -362 12733 -209
rect 13181 -362 13197 -195
rect 10116 -382 10317 -372
rect 12715 -377 13197 -362
rect 10116 -534 10317 -524
rect 5213 -1109 9745 -1059
rect 9819 -586 10116 -536
rect 5012 -1130 5213 -1120
rect 9495 -1180 9768 -1179
rect 3481 -1192 9768 -1180
rect 3481 -1421 9505 -1192
rect 3481 -1422 7466 -1421
rect 3481 -1560 4621 -1422
rect 4768 -1560 5199 -1422
rect 5346 -1424 6835 -1422
rect 5346 -1560 5760 -1424
rect 3481 -1562 5760 -1560
rect 5907 -1560 6835 -1424
rect 6982 -1559 7466 -1422
rect 8289 -1559 9505 -1421
rect 6982 -1560 9505 -1559
rect 5907 -1562 9505 -1560
rect 3481 -1565 9505 -1562
rect 9756 -1565 9768 -1192
rect 3481 -1577 9768 -1565
rect 3481 -1578 9715 -1577
rect 3481 -1874 4114 -1578
rect 6690 -1643 6891 -1633
rect 9819 -1650 9869 -586
rect 10317 -586 10375 -536
rect 10116 -609 10317 -599
rect 6891 -1700 9869 -1650
rect 6690 -1718 6891 -1708
rect 3481 -1886 11682 -1874
rect 3481 -1887 10357 -1886
rect 3481 -2018 9509 -1887
rect 2460 -2023 9509 -2018
rect 2460 -2144 4622 -2023
rect 8372 -2144 9509 -2023
rect 2460 -2222 9509 -2144
rect 9963 -2222 10357 -1887
rect 2460 -2224 10357 -2222
rect 11571 -2224 11682 -1886
rect 2460 -2415 11682 -2224
use sky130_fd_pr__diode_pd2nw_05v5_K4SERG  D1
timestamp 1698886478
transform 1 0 3817 0 1 -1177
box -321 -321 321 321
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D2
timestamp 1698886478
transform 1 0 3679 0 1 -410
box -183 -183 183 183
use level_shifter  level_shifter_0
timestamp 1698887706
transform -1 0 12772 0 1 342
box -422 -2464 2656 76
use level_shifter  level_shifter_1
timestamp 1698887706
transform -1 0 12772 0 -1 470
box -422 -2464 2656 76
use sky130_fd_pr__pfet_01v8_LGS3BL  sky130_fd_pr__pfet_01v8_LGS3BL_0
timestamp 1698716925
transform 0 1 13002 -1 0 643
box -211 -284 211 284
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM1
timestamp 1698886478
transform 1 0 5950 0 1 -1190
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM2
timestamp 1698886478
transform 1 0 6174 0 1 -367
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM3
timestamp 1698886478
transform 1 0 6790 0 1 -367
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM4
timestamp 1698886478
transform 1 0 7062 0 1 -1190
box -278 -300 278 300
use sky130_fd_pr__nfet_01v8_L9WNCD  XM5
timestamp 1699029959
transform 0 1 12859 -1 0 169
box -211 -229 211 229
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM9
timestamp 1698886478
transform 1 0 7406 0 1 -367
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM10
timestamp 1698886478
transform 1 0 7618 0 1 -1190
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM11
timestamp 1698886478
transform 1 0 8022 0 1 -367
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM12
timestamp 1698886478
transform 1 0 8174 0 1 -1190
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM13
timestamp 1698886478
transform 1 0 7062 0 1 -1790
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM14
timestamp 1698886478
transform 1 0 8638 0 1 -367
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM21
timestamp 1698886478
transform 1 0 4838 0 1 -1790
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM22
timestamp 1698886478
transform 1 0 4942 0 1 -367
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM23
timestamp 1698886478
transform 1 0 4838 0 1 -1190
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM24
timestamp 1698886478
transform 1 0 5558 0 1 -367
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM29
timestamp 1698886478
transform 1 0 5950 0 1 -1790
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM30
timestamp 1698886478
transform 1 0 5394 0 1 -1790
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM31
timestamp 1698886478
transform 1 0 7618 0 1 -1790
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM33
timestamp 1698886478
transform 1 0 6506 0 1 -1790
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM34
timestamp 1698886478
transform 1 0 4326 0 1 -367
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM36
timestamp 1698886478
transform 1 0 5394 0 1 -1190
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM39
timestamp 1698886478
transform 1 0 8174 0 1 -1790
box -278 -300 278 300
use sky130_fd_pr__res_xhigh_po_0p35_CWLS5Y  XR1
timestamp 1698886478
transform 1 0 3746 0 1 1544
box -948 -1382 948 1382
use sky130_fd_pr__res_xhigh_po_0p35_7RFGLT  XR2
timestamp 1698886478
transform 1 0 3156 0 1 -1012
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_4FEQLC  XR3
timestamp 1698886478
transform 1 0 7161 0 1 1542
box -2193 -1382 2193 1382
use sky130_fd_pr__res_xhigh_po_0p35_ENTFM9  XR4
timestamp 1699029959
transform 1 0 9281 0 1 -1015
box -284 -1082 284 1082
use sky130_fd_pr__res_xhigh_po_0p35_KNBXRF  XR5
timestamp 1698886478
transform 1 0 9801 0 1 1342
box -201 -1582 201 1582
<< labels >>
flabel metal2 2460 -2415 2662 -790 0 FreeSans 256 0 0 0 avss
port 3 nsew
flabel metal1 2460 -722 2660 -522 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 2460 1016 2660 1216 0 FreeSans 256 0 0 0 in
port 0 nsew
flabel metal2 2460 1587 2585 3215 0 FreeSans 256 0 0 0 avdd
port 2 nsew
flabel metal2 13186 418 13386 1190 0 FreeSans 256 0 0 0 dvdd
port 4 nsew
flabel metal1 13168 -2348 13364 -1384 0 FreeSans 256 0 0 0 dvss
port 5 nsew
flabel metal1 13164 -962 13364 -762 0 FreeSans 256 0 0 0 ena
port 6 nsew
flabel metal1 13164 1574 13364 1774 0 FreeSans 256 0 0 0 stdby
port 8 nsew
flabel metal1 13164 88 13364 288 0 FreeSans 256 0 0 0 dout
port 7 nsew
<< end >>
