magic
tech sky130A
magscale 1 2
timestamp 1699029959
<< pwell >>
rect -284 -1082 284 1082
<< psubdiff >>
rect -248 1012 -152 1046
rect 152 1012 248 1046
rect -248 950 -214 1012
rect 214 950 248 1012
rect -248 -1012 -214 -950
rect 214 -1012 248 -950
rect -248 -1046 -152 -1012
rect 152 -1046 248 -1012
<< psubdiffcont >>
rect -152 1012 152 1046
rect -248 -950 -214 950
rect 214 -950 248 950
rect -152 -1046 152 -1012
<< xpolycontact >>
rect -118 484 -48 916
rect -118 -916 -48 -484
rect 48 484 118 916
rect 48 -916 118 -484
<< xpolyres >>
rect -118 -484 -48 484
rect 48 -484 118 484
<< locali >>
rect -248 1012 -152 1046
rect 152 1012 248 1046
rect -248 950 -214 1012
rect 214 950 248 1012
rect -248 -1012 -214 -950
rect 214 -1012 248 -950
rect -248 -1046 -152 -1012
rect 152 -1046 248 -1012
<< viali >>
rect -102 501 -64 898
rect 64 501 102 898
rect -102 -898 -64 -501
rect 64 -898 102 -501
<< metal1 >>
rect -108 898 -58 910
rect -108 501 -102 898
rect -64 501 -58 898
rect -108 489 -58 501
rect 58 898 108 910
rect 58 501 64 898
rect 102 501 108 898
rect 58 489 108 501
rect -108 -501 -58 -489
rect -108 -898 -102 -501
rect -64 -898 -58 -501
rect -108 -910 -58 -898
rect 58 -501 108 -489
rect 58 -898 64 -501
rect 102 -898 108 -501
rect 58 -910 108 -898
<< properties >>
string FIXED_BBOX -231 -1029 231 1029
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 5.0 m 1 nx 2 wmin 0.350 lmin 0.50 rho 2000 val 29.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
